module print_table(
    input wire clk,           // ��ȷ��ʱ��Ƶ�ʣ�Ĭ�ϰ� 100MHz ��д
    input wire rst_n,
    input wire start,         // �ⲿ��������
    // UART TX �ӿ�
    input wire uart_tx_busy,
    output reg uart_tx_en,
    output reg [7:0] uart_tx_data,
    // ��������
    input wire [49:0] info_table,
    input wire [7:0] cnt,     
    output reg busy,
    output reg done,
    output reg [3:0] current_state
);

    // --- ASCII ���� ---
    localparam [7:0] ASCII_STAR  = 8'h2A, ASCII_SPACE = 8'h20,
                     ASCII_0     = 8'h30, ASCII_CR    = 8'h0D, ASCII_LF = 8'h0A;

    // --- ״̬������ ---
    localparam S_IDLE        = 4'd0,
               S_PREPARE     = 4'd1,
               S_SET_DATA    = 4'd2,
               S_SEND_TRIG   = 4'd3,
               S_WAIT_START  = 4'd4, // �ȴ� busy ����
               S_WAIT_DONE   = 4'd5, // �ȴ� busy ����
               S_COOL_DOWN   = 4'd6, // ǿ����ȴ����ֹ�������絼������
               S_DONE        = 4'd7;

    reg [3:0] state, next_state;
    reg [5:0] step_cnt; 
    reg [4:0] cell_idx; 
    reg [2:0] row, col; 
    reg [7:0] t_tens, t_ones;
    reg [1:0] cur_cell_val;
    reg [19:0] cool_cnt; // ��ȴ������

    // ��ȴʱ�䳣����100,000 �������� 100MHz �µ��� 1ms��ȷ�������߾��Կ���
    localparam COOL_TIME = 20'd100_000; 

    wire [4:0] cur_place = (col - 3'd1) * 3'd5 + (row - 3'd1);

    // --- ��һ�Σ�ʱ���߼� ---
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) state <= S_IDLE;
        else        state <= next_state;
    end

    // --- �ڶ��Σ�����߼� (��ת����) ---
    always @(*) begin
        next_state = state;
        case (state)
            S_IDLE:       if (start) next_state = S_PREPARE;
            S_PREPARE:    next_state = S_SET_DATA;
            S_SET_DATA:   next_state = S_SEND_TRIG;
            S_SEND_TRIG:  next_state = S_WAIT_START;
            S_WAIT_START: if (uart_tx_busy) next_state = S_WAIT_DONE; // ȷ�����յ�
            S_WAIT_DONE:  if (!uart_tx_busy) next_state = S_COOL_DOWN; // ȷ���ѷ���
            S_COOL_DOWN: begin
                if (cool_cnt >= COOL_TIME) begin
                    if (cell_idx == 5'd25) next_state = S_DONE;
                    else                   next_state = S_SET_DATA;
                end
            end
            S_DONE:       next_state = S_IDLE;
            default:      next_state = S_IDLE;
        endcase
    end

    // --- �����Σ�ʱ���߼� (����·�������) ---
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            uart_tx_en <= 0; uart_tx_data <= 0; busy <= 0; done <= 0;
            step_cnt <= 0; cell_idx <= 0; row <= 1; col <= 1; cool_cnt <= 0;
        end else begin
            case (state)
                S_IDLE: begin
                    busy <= 0; done <= 0; step_cnt <= 0; cell_idx <= 0;
                    row <= 1; col <= 1; cool_cnt <= 0; uart_tx_en <= 0;
                end

                S_PREPARE: begin
                    busy <= 1;
                    t_tens <= cnt / 10;
                    t_ones <= cnt % 10;
                    cur_cell_val <= info_table[49 - (cur_place << 1) -: 2];
                end

                S_SET_DATA: begin
                    cool_cnt <= 0; // ������ȴ����
                    // �����ǰ��ԪcntΪ0�������˵�Ԫ
                    if (cur_cell_val == 2'd0) begin
                        // ֱ��������һ����Ԫ
                        if (col == 3'd5) begin
                            col <= 3'd1;
                            row <= row + 1'b1;
                        end else begin
                            col <= col + 1'b1;
                        end
                        cell_idx <= cell_idx + 1'b1;
                    end else begin
                        case (step_cnt)
                            6'd0:  uart_tx_data <= ASCII_0 + t_tens;
                            6'd1:  uart_tx_data <= ASCII_0 + t_ones;
                            6'd2:  uart_tx_data <= ASCII_SPACE;
                            6'd3:  uart_tx_data <= ASCII_0 + row;
                            6'd4:  uart_tx_data <= ASCII_STAR;
                            6'd5:  uart_tx_data <= ASCII_0 + col;
                            6'd6:  uart_tx_data <= ASCII_STAR;
                            6'd7:  uart_tx_data <= ASCII_0 + cur_cell_val;
                            6'd8:  uart_tx_data <= ASCII_SPACE;
                            6'd9:  uart_tx_data <= ASCII_CR;
                            6'd10: uart_tx_data <= ASCII_LF;
                            default: uart_tx_data <= ASCII_SPACE;
                        endcase
                    end
                end

                S_SEND_TRIG: begin
                    uart_tx_en <= 1'b1;
                end

                S_WAIT_START, S_WAIT_DONE: begin
                    uart_tx_en <= 1'b0;
                end

                S_COOL_DOWN: begin
                    cool_cnt <= cool_cnt + 1'b1;
                    // ����ȴ�ڼ�ĵ�һ�����ڸ�����һ��Ҫ���͵�����
                    if (cool_cnt == 20'd1) begin
                        if (step_cnt < 6'd8) begin
                            step_cnt <= step_cnt + 1'b1;
                        end else if (step_cnt == 6'd8) begin
                            if (col == 3'd5) step_cnt <= 6'd9;
                            else begin
                                step_cnt <= 6'd3; // ��������
                                cell_idx <= cell_idx + 1'b1;
                                col      <= col + 1'b1;
                            end
                        end else if (step_cnt == 6'd9) begin
                            step_cnt <= 6'd10;
                        end else if (step_cnt == 6'd10) begin
                            cell_idx <= cell_idx + 1'b1;
                            if (cell_idx != 5'd24) begin
                                step_cnt <= 6'd3;
                                col <= 3'd1; row <= row + 1'b1;
                            end else begin
                                cell_idx <= 5'd25; // ׼���� DONE
                            end
                        end
                    end
                    // ����ȴ�����ʱ��ǰ������һ�����ݣ���֤ SET_DATA ״̬�����ȶ�
                    if (cool_cnt == COOL_TIME - 1) begin
                        cur_cell_val <= info_table[49 - (cur_place << 1) -: 2];
                    end
                end

                S_DONE: begin
                    done <= 1'b1;
                    busy <= 1'b0;
                end
            endcase
        end
    end

endmodule